bind wb_arbiter arbiter_checker_sva check1(clk, rst, rqst_i, gnt_o);
