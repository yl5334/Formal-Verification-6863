bind wb_arbiter arbiter_checker_ovl check0(clk, rst, rqst_i, gnt_o);
